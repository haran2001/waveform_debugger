//--------------DESCRIPTION--------------
// This is a testbench for the FIFO module.
// The testbench generates random data and writes it to the FIFO, 
// then reads it back and compares the results.
//---------------------------------------

`timescale 1ns/1ps

module FIFO_tb();

    parameter DSIZE = 8; // Data bus size
    parameter ASIZE = 3; // Address bus size
    parameter DEPTH = 1 << ASIZE; // Depth of the FIFO memory

    reg [DSIZE-1:0] wdata;   // Input data
    wire [DSIZE-1:0] rdata;  // Output data
    wire wfull, rempty;      // Write full and read empty signals
    reg winc, rinc, wclk, rclk, wrst_n, rrst_n; // Write and read signals

    FIFO #(DSIZE, ASIZE) fifo (
        .rdata(rdata), 
        .wdata(wdata),
        .wfull(wfull),
        .rempty(rempty),
        .winc(winc), 
        .rinc(rinc), 
        .wclk(wclk), 
        .rclk(rclk), 
        .wrst_n(wrst_n), 
        .rrst_n(rrst_n)
    );

    integer i=0;
    integer seed = 1;

    // Read and write clock in loop
    always #5 wclk = ~wclk;    // faster writing
    always #10 rclk = ~rclk;   // slower reading
    
    initial begin
        // Initialize all signals
        wclk = 0;
        rclk = 0;
        wrst_n = 1;     // Active low reset
        rrst_n = 1;     // Active low reset
        winc = 0;
        rinc = 0;
        wdata = 0;

        // Reset the FIFO
        #40 wrst_n = 0; rrst_n = 0;
        #40 wrst_n = 1; rrst_n = 1;

        // TEST CASE 1: Write data and read it back
        rinc = 1;
        for (i = 0; i < 10; i = i + 1) begin
            wdata = $random(seed) % 256;
            winc = 1;
            #10;
            winc = 0;
            #10;
        end

        // TEST CASE 2: Write data to make FIFO full and try to write more data
        rinc = 0;
        winc = 1;
        for (i = 0; i < DEPTH + 3; i = i + 1) begin
            wdata = $random(seed) % 256;
            #10;
        end

        // Add after TEST CASE 2 (around line 70), before TEST CASE 3:

        // Try one more write while full - should be blocked
        wdata = 8'hFF;
        winc = 1;
        #10;
        winc = 0;
        #10;

        // Verify wfull still asserted (no overflow occurred)
        if (!wfull) begin
            $display("FAIL: wfull deasserted after write attempt at t=%0t. Possible overflow.", $time);
            $fatal;
        end

        // TEST CASE 3: Read data from empty FIFO and try to read more data
        winc = 0;
        rinc = 1;
        for (i = 0; i < DEPTH + 3; i = i + 1) begin
            #20;
        end

        // TEST CASE 4: Strict wfull timing verification
        $display("\n--- TEST CASE 4: wfull timing verification ---");

        // Reset FIFO first
        wrst_n = 0; rrst_n = 0;
        #40;
        wrst_n = 1; rrst_n = 1;
        #40;

        rinc = 0;
        winc = 0;

        // Verify wfull is 0 when empty
        if (wfull) begin
            $display("FAIL: wfull=1 after reset at t=%0t. Expected wfull=0 for empty FIFO", $time);
            $fatal;
        end

        // Fill FIFO one entry at a time, checking wfull each time
        for (i = 0; i < DEPTH; i = i + 1) begin
            // wfull should be 0 before FIFO is full
            if (wfull) begin
                $display("FAIL: wfull asserted too early at t=%0t after %0d writes. Expected wfull=0 until %0d writes.", 
                        $time, i, DEPTH);
                $fatal;
            end
            
            wdata = i; // Use index as data for easy tracking
            winc = 1;
            #10;
            winc = 0;
            #10;
        end

        // Now FIFO has exactly DEPTH entries - wfull MUST be 1
        #20; // Allow for synchronizer delay
        if (!wfull) begin
            $display("FAIL: wfull not asserted at t=%0t after %0d writes. wfull=%b, expected=1", 
                    $time, DEPTH, wfull);
            $fatal;
        end

        $display("PASS: wfull correctly asserted after exactly %0d writes at t=%0t", DEPTH, $time);


        $finish;
    end

endmodule

//----------------------------EXPLANATION-----------------------------------------------
// The testbench for the FIFO module generates random data and writes it to the FIFO,
// then reads it back and compares the results. The testbench includes three test cases:
// 1. Write data and read it back.
// 2. Write data to make the FIFO full and try to write more data.
// 3. Read data from an empty FIFO and try to read more data. The testbench uses
// clock signals for writing and reading, and includes reset signals to initialize
// the FIFO. The testbench finishes after running the test cases.
//--------------------------------------------------------------------------------------
